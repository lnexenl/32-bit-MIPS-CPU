`timescale 1ns/1ps

module ROM (addr,data);
input [30:0] addr;
output [31:0] data;

localparam ROM_SIZE = 150;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data=(addr < (ROM_SIZE << 2))?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin
ROMDATA[0] <= 32'h8000003;
ROMDATA[1] <= 32'h800002d;
ROMDATA[2] <= 32'h800002c;
ROMDATA[3] <= 32'h3c084000;
ROMDATA[4] <= 32'h8d090020;
ROMDATA[5] <= 32'h31290002;
ROMDATA[6] <= 32'h1120fffd;
ROMDATA[7] <= 32'h8d10001c;
ROMDATA[8] <= 32'h8d090020;
ROMDATA[9] <= 32'h31290002;
ROMDATA[10] <= 32'h1120fffd;
ROMDATA[11] <= 32'h8d11001c;
ROMDATA[12] <= 32'had000008;
ROMDATA[13] <= 32'h2009fc18;
ROMDATA[14] <= 32'had090000;
ROMDATA[15] <= 32'had090004;
ROMDATA[16] <= 32'h20090003;
ROMDATA[17] <= 32'had090008;
ROMDATA[18] <= 32'h10b020;
ROMDATA[19] <= 32'h11b820;
ROMDATA[20] <= 32'h200f0001;
ROMDATA[21] <= 32'h800001c;
ROMDATA[22] <= 32'h11000001;
ROMDATA[23] <= 32'h11200002;
ROMDATA[24] <= 32'h108042;
ROMDATA[25] <= 32'h800001c;
ROMDATA[26] <= 32'h118842;
ROMDATA[27] <= 32'h800001c;
ROMDATA[28] <= 32'h32080001;
ROMDATA[29] <= 32'h32290001;
ROMDATA[30] <= 32'h1095020;
ROMDATA[31] <= 32'h114ffff6;
ROMDATA[32] <= 32'h12110008;
ROMDATA[33] <= 32'h211402a;
ROMDATA[34] <= 32'h11000003;
ROMDATA[35] <= 32'h2308822;
ROMDATA[36] <= 32'h12110004;
ROMDATA[37] <= 32'h800001c;
ROMDATA[38] <= 32'h2118022;
ROMDATA[39] <= 32'h12110001;
ROMDATA[40] <= 32'h800001c;
ROMDATA[41] <= 32'h3c124000;
ROMDATA[42] <= 32'hae500018;
ROMDATA[43] <= 32'h800002b;
ROMDATA[44] <= 32'h3600008;
ROMDATA[45] <= 32'hae50000c;
ROMDATA[46] <= 32'h8e530008;
ROMDATA[47] <= 32'h2014fff9;
ROMDATA[48] <= 32'h2749824;
ROMDATA[49] <= 32'hae530008;
ROMDATA[50] <= 32'h22520014;
ROMDATA[51] <= 32'h8e530000;
ROMDATA[52] <= 32'h32730f00;
ROMDATA[53] <= 32'h20140100;
ROMDATA[54] <= 32'h10140007;
ROMDATA[55] <= 32'h1274000a;
ROMDATA[56] <= 32'h14a040;
ROMDATA[57] <= 32'h1274000d;
ROMDATA[58] <= 32'h14a040;
ROMDATA[59] <= 32'h1274000f;
ROMDATA[60] <= 32'h14a040;
ROMDATA[61] <= 32'h12740000;
ROMDATA[62] <= 32'h20140100;
ROMDATA[63] <= 32'h32cc000f;
ROMDATA[64] <= 32'hc000050;
ROMDATA[65] <= 32'h800008e;
ROMDATA[66] <= 32'h14a040;
ROMDATA[67] <= 32'h32cc00f0;
ROMDATA[68] <= 32'hc6102;
ROMDATA[69] <= 32'hc000050;
ROMDATA[70] <= 32'h800008e;
ROMDATA[71] <= 32'h14a040;
ROMDATA[72] <= 32'h32ec000f;
ROMDATA[73] <= 32'hc000050;
ROMDATA[74] <= 32'h800008e;
ROMDATA[75] <= 32'h14a040;
ROMDATA[76] <= 32'h32ec00f0;
ROMDATA[77] <= 32'hc6102;
ROMDATA[78] <= 32'hc000050;
ROMDATA[79] <= 32'h800008e;
ROMDATA[80] <= 32'h9820;
ROMDATA[81] <= 32'h1193001e;
ROMDATA[82] <= 32'h22730001;
ROMDATA[83] <= 32'h1193001e;
ROMDATA[84] <= 32'h22730001;
ROMDATA[85] <= 32'h1193001e;
ROMDATA[86] <= 32'h22730001;
ROMDATA[87] <= 32'h1193001e;
ROMDATA[88] <= 32'h22730001;
ROMDATA[89] <= 32'h1193001e;
ROMDATA[90] <= 32'h22730001;
ROMDATA[91] <= 32'h1193001e;
ROMDATA[92] <= 32'h22730001;
ROMDATA[93] <= 32'h1193001e;
ROMDATA[94] <= 32'h22730001;
ROMDATA[95] <= 32'h1193001e;
ROMDATA[96] <= 32'h22730001;
ROMDATA[97] <= 32'h1193001e;
ROMDATA[98] <= 32'h22730001;
ROMDATA[99] <= 32'h1193001e;
ROMDATA[100] <= 32'h22730001;
ROMDATA[101] <= 32'h1193001e;
ROMDATA[102] <= 32'h22730001;
ROMDATA[103] <= 32'h1193001e;
ROMDATA[104] <= 32'h22730001;
ROMDATA[105] <= 32'h1193001e;
ROMDATA[106] <= 32'h22730001;
ROMDATA[107] <= 32'h1193001e;
ROMDATA[108] <= 32'h22730001;
ROMDATA[109] <= 32'h1193001e;
ROMDATA[110] <= 32'h200c0071;
ROMDATA[111] <= 32'h3e00008;
ROMDATA[112] <= 32'h200c003f;
ROMDATA[113] <= 32'h3e00008;
ROMDATA[114] <= 32'h200c0006;
ROMDATA[115] <= 32'h3e00008;
ROMDATA[116] <= 32'h200c005b;
ROMDATA[117] <= 32'h3e00008;
ROMDATA[118] <= 32'h200c004f;
ROMDATA[119] <= 32'h3e00008;
ROMDATA[120] <= 32'h200c0066;
ROMDATA[121] <= 32'h3e00008;
ROMDATA[122] <= 32'h200c006d;
ROMDATA[123] <= 32'h3e00008;
ROMDATA[124] <= 32'h200c007d;
ROMDATA[125] <= 32'h3e00008;
ROMDATA[126] <= 32'h200c0007;
ROMDATA[127] <= 32'h3e00008;
ROMDATA[128] <= 32'h200c007f;
ROMDATA[129] <= 32'h3e00008;
ROMDATA[130] <= 32'h200c006f;
ROMDATA[131] <= 32'h3e00008;
ROMDATA[132] <= 32'h200c0077;
ROMDATA[133] <= 32'h3e00008;
ROMDATA[134] <= 32'h200c007c;
ROMDATA[135] <= 32'h3e00008;
ROMDATA[136] <= 32'h200c0039;
ROMDATA[137] <= 32'h3e00008;
ROMDATA[138] <= 32'h200c005e;
ROMDATA[139] <= 32'h3e00008;
ROMDATA[140] <= 32'h200c0079;
ROMDATA[141] <= 32'h3e00008;
ROMDATA[142] <= 32'h1946020;
ROMDATA[143] <= 32'hae4c0000;
ROMDATA[144] <= 32'h2252fff4;
ROMDATA[145] <= 32'h8e530000;
ROMDATA[146] <= 32'h20140002;
ROMDATA[147] <= 32'h2749825;
ROMDATA[148] <= 32'hae530000;
ROMDATA[149] <= 32'h3400008;

end
endmodule
