module ALU(A,B,Z,Sign,ALUFun);
input [31:0] A;
input [31:0] B;
input [5:0] ALUFun;
input Sign;
output reg[31:0] Z;
wire [31:0] Z1,Z2;
wire V=1'b0,V1=1'b0,V2=1'b0;
wire N=1'b0,N1=1'b0,N2=1'b0;
wire 
ADDER(A,B,Sign,Z1,V1,N1)
ADDER(A,~B,Sign,Z2,V2,N2)
	always @(*)
		case (ALUFun)
// compute
			6'b000000:
			begin
				Z <= Z1;
				V <= V1;
				N <= N1;
			end
			6'b000001:
			begin
			  Z <= Z2;
			  V <= V2;
			  N <= N2;
			end 
// logic
			6'b011000: Z <= A & B;
			6'b011110: Z <= A | B;
			6'b010110: Z <= A ^ B;
			6'b010001: Z <=~(A|B);
			6'b011010: Z <= A    ;
//changeposition
			6'b100000: 
			begin
			  if(A[0]) B << 1;
			  if(A[1]) B << 2;
			  if(A[2]) B << 4;
			  if(A[3]) B << 8;
			  if(A[4]) B << 16;
			end 
			6'b100001:
			begin
			  if(A[0]) B >> 1;
			  if(A[1]) B >> 2;
			  if(A[2]) B >> 4;
			  if(A[3]) B >> 8;
			  if(A[4]) B >> 16;
			end
			6'b100011:
			begin
			  BB[31:0] <= B;
			  BB[32] <= BB[31];
			  if(A[0]) BB >> 1;
			  if(A[1]) BB >> 2;
			  if(A[2]) BB >> 4;
			  if(A[3]) BB >> 8;
			  if(A[4]) BB >> 16;
			  B <= BB[31:0];
			end 
//corleration
			6'b110011:
			begin
			  	Z <= (N2==1'b1)?32'b0000_0000_0000_0000_0000_0000_0000_0001:8'h00000000;
			end 
			6'b110001: Z <= (N2!=1'b1)?32'b0000_0000_0000_0000_0000_0000_0000_0001:8'h00000000;
			6'b110101: Z <= (V2==1'b1)?32'b0000_0000_0000_0000_0000_0000_0000_0001:8'h00000000;
			6'b111101: Z <= ((Sign==1'b1&&A[31]==1'b1)||A==8'h00000000||A==32'b1000_0000_0000_0000_0000_0000_0000_0000)?32'b0000_0000_0000_0000_0000_0000_0000_0001:8'h00000000;
			6'b111011: Z <= (Sign==1'b1&&A[31]==1'b1)?32'b0000_0000_0000_0000_0000_0000_0000_0001:8'h00000000;
			6'b111111: Z <= (((Sign==1'b1&&A[31]==1'b0)||(Sign==1'b0))&&(A!=8'h00000000))?32'b0000_0000_0000_0000_0000_0000_0000_0001:8'h00000000;
			default: Z <= 32'h00000000;
		endcase

endmodule