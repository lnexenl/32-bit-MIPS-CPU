`timescale 1ns/1ps

module ROM (addr,data);
input [30:0] addr;
output [31:0] data;

localparam ROM_SIZE = 137;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data=(addr < ROM_SIZE)?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin
		ROMDATA[0] <= 32'h800000c;
ROMDATA[1] <= 32'h8000022;
ROMDATA[2] <= 32'h8000021;
ROMDATA[3] <= 32'h211ffc18;
ROMDATA[4] <= 32'h3c084009;
ROMDATA[5] <= 32'had090000;
ROMDATA[6] <= 32'h21080004;
ROMDATA[7] <= 32'had090000;
ROMDATA[8] <= 32'h21080004;
ROMDATA[9] <= 32'had000000;
ROMDATA[10] <= 32'h22000002;
ROMDATA[11] <= 32'h22200004;
ROMDATA[12] <= 32'h21e00001;
ROMDATA[13] <= 32'h8000014;
ROMDATA[14] <= 32'h10fffffe;
ROMDATA[15] <= 32'h111ffffd;
ROMDATA[16] <= 32'h108042;
ROMDATA[17] <= 32'h8000014;
ROMDATA[18] <= 32'h118842;
ROMDATA[19] <= 32'h8000014;
ROMDATA[20] <= 32'h31100001;
ROMDATA[21] <= 32'h31310001;
ROMDATA[22] <= 32'h1095020;
ROMDATA[23] <= 32'h114f0009;
ROMDATA[24] <= 32'h1210fff7;
ROMDATA[25] <= 32'h211402a;
ROMDATA[26] <= 32'h10fffffc;
ROMDATA[27] <= 32'h2308822;
ROMDATA[28] <= 32'h1210fffb;
ROMDATA[29] <= 32'h8000014;
ROMDATA[30] <= 32'h2118022;
ROMDATA[31] <= 32'h1210fffe;
ROMDATA[32] <= 32'h8000014;
ROMDATA[33] <= 32'h3600008;
ROMDATA[34] <= 32'h3c124009;
ROMDATA[35] <= 32'h22520008;
ROMDATA[36] <= 32'h8e530000;
ROMDATA[37] <= 32'h227ffff9;
ROMDATA[38] <= 32'h2749824;
ROMDATA[39] <= 32'hae530000;
ROMDATA[40] <= 32'h2252000c;
ROMDATA[41] <= 32'h8e530000;
ROMDATA[42] <= 32'h32730f00;
ROMDATA[43] <= 32'h22800100;
ROMDATA[44] <= 32'h1273ffef;
ROMDATA[45] <= 32'h14a040;
ROMDATA[46] <= 32'h1273ffec;
ROMDATA[47] <= 32'h14a040;
ROMDATA[48] <= 32'h1273ffe9;
ROMDATA[49] <= 32'h14a040;
ROMDATA[50] <= 32'h1273fffc;
ROMDATA[51] <= 32'h14a0c2;
ROMDATA[52] <= 32'h3190000f;
ROMDATA[53] <= 32'hc00004c;
ROMDATA[54] <= 32'h800008b;
ROMDATA[55] <= 32'h14a040;
ROMDATA[56] <= 32'h319000f0;
ROMDATA[57] <= 32'hc00004c;
ROMDATA[58] <= 32'h800008b;
ROMDATA[59] <= 32'h14a040;
ROMDATA[60] <= 32'h3191000f;
ROMDATA[61] <= 32'hc00004c;
ROMDATA[62] <= 32'h800008b;
ROMDATA[63] <= 32'h14a040;
ROMDATA[64] <= 32'h319100f0;
ROMDATA[65] <= 32'hc00004c;
ROMDATA[66] <= 32'h800008b;
ROMDATA[67] <= 32'h9820;
ROMDATA[68] <= 32'h1192ffd7;
ROMDATA[69] <= 32'h22730001;
ROMDATA[70] <= 32'h1192ffd7;
ROMDATA[71] <= 32'h22730001;
ROMDATA[72] <= 32'h1192ffd7;
ROMDATA[73] <= 32'h22730001;
ROMDATA[74] <= 32'h1192ffd7;
ROMDATA[75] <= 32'h22730001;
ROMDATA[76] <= 32'h1192ffd7;
ROMDATA[77] <= 32'h22730001;
ROMDATA[78] <= 32'h1192ffd7;
ROMDATA[79] <= 32'h22730001;
ROMDATA[80] <= 32'h1192ffd7;
ROMDATA[81] <= 32'h22730001;
ROMDATA[82] <= 32'h1192ffd7;
ROMDATA[83] <= 32'h22730001;
ROMDATA[84] <= 32'h1192ffd7;
ROMDATA[85] <= 32'h22730001;
ROMDATA[86] <= 32'h1192ffd7;
ROMDATA[87] <= 32'h22730001;
ROMDATA[88] <= 32'h1192ffd7;
ROMDATA[89] <= 32'h22730001;
ROMDATA[90] <= 32'h1192ffd7;
ROMDATA[91] <= 32'h22730001;
ROMDATA[92] <= 32'h1192ffd7;
ROMDATA[93] <= 32'h22730001;
ROMDATA[94] <= 32'h1192ffd7;
ROMDATA[95] <= 32'h22730001;
ROMDATA[96] <= 32'h1192ffd7;
ROMDATA[97] <= 32'h21800071;
ROMDATA[98] <= 32'h3e00008;
ROMDATA[99] <= 32'h2180003f;
ROMDATA[100] <= 32'h3e00008;
ROMDATA[101] <= 32'h21800006;
ROMDATA[102] <= 32'h3e00008;
ROMDATA[103] <= 32'h2180005b;
ROMDATA[104] <= 32'h3e00008;
ROMDATA[105] <= 32'h2180004f;
ROMDATA[106] <= 32'h3e00008;
ROMDATA[107] <= 32'h21800066;
ROMDATA[108] <= 32'h3e00008;
ROMDATA[109] <= 32'h2180006d;
ROMDATA[110] <= 32'h3e00008;
ROMDATA[111] <= 32'h2180007d;
ROMDATA[112] <= 32'h3e00008;
ROMDATA[113] <= 32'h21800007;
ROMDATA[114] <= 32'h3e00008;
ROMDATA[115] <= 32'h2180007f;
ROMDATA[116] <= 32'h3e00008;
ROMDATA[117] <= 32'h2180006f;
ROMDATA[118] <= 32'h3e00008;
ROMDATA[119] <= 32'h21800077;
ROMDATA[120] <= 32'h3e00008;
ROMDATA[121] <= 32'h2180007c;
ROMDATA[122] <= 32'h3e00008;
ROMDATA[123] <= 32'h21800039;
ROMDATA[124] <= 32'h3e00008;
ROMDATA[125] <= 32'h2180005e;
ROMDATA[126] <= 32'h3e00008;
ROMDATA[127] <= 32'h21800079;
ROMDATA[128] <= 32'h3e00008;
ROMDATA[129] <= 32'h1946020;
ROMDATA[130] <= 32'hae4c0000;
ROMDATA[131] <= 32'h2251fff4;
ROMDATA[132] <= 32'h8e530000;
ROMDATA[133] <= 32'h22800002;
ROMDATA[134] <= 32'h2749825;
ROMDATA[135] <= 32'hae530000;
ROMDATA[136] <= 32'h3400008;
end
endmodule
